typedef enum logic [2:0] {
    ADD,
    SUB,
    MUL,
    DIV,
    AND,
    OR,
    XOR
} alu_functions_e;
module alu ();
endmodule
