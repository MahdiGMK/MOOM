module multiplier ();

endmodule
