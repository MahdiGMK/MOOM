module alu ();
  adder #(.NBIT(10)) test_adder ();
endmodule
