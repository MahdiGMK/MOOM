module test ();
endmodule
// verilator lint_off DECLFILENAME
